/************************************************************************
Avalon-MM Interface for AES Decryption IP Core

Dong Kai Wang, Fall 2017

For use with ECE 385 Experiment 9
University of Illinois ECE Department

Register Map:

 0-3 : 4x 32bit AES Key
 4-7 : 4x 32bit AES Encrypted Message
 8-11: 4x 32bit AES Decrypted Message
   12: Not Used
	13: Not Used
   14: 32bit Start Register
   15: 32bit Done Register

************************************************************************/

module avalon_aes_interface (
	// Avalon Clock Input
	input logic CLK,
	
	// Avalon Reset Input
	input logic RESET,
	
	// Avalon-MM Slave Signals
	input  logic AVL_READ,					// Avalon-MM Read
	input  logic AVL_WRITE,					// Avalon-MM Write
	input  logic AVL_CS,						// Avalon-MM Chip Select
	input  logic [3:0] AVL_BYTE_EN,		// Avalon-MM Byte Enable
	input  logic [3:0] AVL_ADDR,			// Avalon-MM Address
	input  logic [31:0] AVL_WRITEDATA,	// Avalon-MM Write Data
	output logic [31:0] AVL_READDATA,	// Avalon-MM Read Data
	
	// Exported Conduit
	output logic [31:0] EXPORT_DATA		// Exported Conduit Signal to LEDs
);
	
	logic[31:0] regs[16];
	logic[31:0] regs2[4];
	logic done;
		AES Decryption_Logic(.CLK(CLK),.RESET(RESET),.AES_START(regs[14][0]),
						.AES_DONE(done),.AES_KEY({regs[0][31:0],regs[1][31:0],regs[2][31:0],regs[3][31:0]}),
						.AES_MSG_ENC({regs[4][31:0],regs[5][31:0],regs[6][31:0],regs[7][31:0]}),
						.AES_MSG_DEC({regs2[0],regs2[1],regs2[2],regs2[3]})
);

			always_ff @ (posedge CLK)
				begin
				if(RESET)
					begin
						for(int i=0;i<16;i++)
						begin 
							regs[i] <= 32'b0;
						end
					end
					if(AVL_WRITE == 1'b1 && AVL_CS == 1'b1)
						begin
						case (AVL_BYTE_EN)
						4'b1100:begin regs[AVL_ADDR][31:16] <= AVL_WRITEDATA[31:16]; end
						4'b0011:begin regs[AVL_ADDR][15:0] <= AVL_WRITEDATA[15:0]; end
						4'b1000:begin regs[AVL_ADDR][31:24] <= AVL_WRITEDATA[31:24];end
						4'b0100:begin regs[AVL_ADDR][23:16] <= AVL_WRITEDATA[23:16];end
						4'b0010:begin regs[AVL_ADDR][15:7] <= AVL_WRITEDATA[15:7];end 
						4'b0001:begin regs[AVL_ADDR][7:0] <= AVL_WRITEDATA[7:0]; end
						default:begin regs[AVL_ADDR] <= AVL_WRITEDATA;end
						endcase
						end
					if(done)
					begin
					regs[8][31:0] <= regs2[0];
					regs[9][31:0] <= regs2[1];
					regs[10][31:0] <= regs2[2];
					regs[11][31:0] <= regs2[3];
					regs[15][0] <= done;
					end
				end
				
				always_comb
				begin
					if(AVL_READ == 1'b1 && AVL_CS == 1'b1)
					begin
						AVL_READDATA = regs[AVL_ADDR];
					end
					else
					begin 
						AVL_READDATA = 32'hXXXXXXXX;
					end
				end
			assign EXPORT_DATA[31:16] = regs[4][31:16];
			assign EXPORT_DATA[15:0] = regs[7][15:0];

endmodule
